module Timer (
	state,
	sig_Full,
	sig_Temperature,
	sig_Completed
	);
	
	input [2:0] state;
	output sig_Full;
	output sig_Temperature;
	output sig_Completed;
	




endmodule
